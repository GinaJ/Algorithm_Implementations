library ieee;
use ieee.std_logic_1164.all;

package myTypes is
    
    --Define size of a single number-->number of bit 
    constant NBIT : natural := 16;    
    
    --Define size of the CUBE (size of i, j, k)
    constant i_size :=3;
    constant j_size :=3;
    constant k_size :=3;
    
    end myTypes;